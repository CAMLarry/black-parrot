// Top level TAGE

//

// controller

// incrementer

// branch address

// index tag gen

// bimodal table

// tage table x4

// 4x comparators

// update predictor

// update history

// 