module local_history_table ();

