// branch